library verilog;
use verilog.vl_types.all;
entity ALUtest is
end ALUtest;
