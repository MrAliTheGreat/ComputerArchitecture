library verilog;
use verilog.vl_types.all;
entity TestBench_DataPath is
end TestBench_DataPath;
