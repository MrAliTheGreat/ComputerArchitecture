library verilog;
use verilog.vl_types.all;
entity TestBench_12_bit is
end TestBench_12_bit;
