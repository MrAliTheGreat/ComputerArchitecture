library verilog;
use verilog.vl_types.all;
entity DATAPATH is
    port(
        clk             : in     vl_logic
    );
end DATAPATH;
