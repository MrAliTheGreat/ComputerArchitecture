library verilog;
use verilog.vl_types.all;
entity PDP_8 is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end PDP_8;
