library verilog;
use verilog.vl_types.all;
entity tb_datapath is
end tb_datapath;
