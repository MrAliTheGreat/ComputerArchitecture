`timescale 1ns/1ns
module Adder_6_bit(input [5:0] y , input[5:0] p , output [5:0] Q);
  assign Q = y + p;

endmodule
