library verilog;
use verilog.vl_types.all;
entity TestBench_Controller is
end TestBench_Controller;
