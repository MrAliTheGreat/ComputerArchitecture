`timescale 1ns/1ns
module tb_datapath ();
 
  reg clk = 1'b1;
 
  DATAPATH uut (clk);
  
  initial begin
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
    #100 clk = ~clk;#100 clk = ~clk;
  end
endmodule

